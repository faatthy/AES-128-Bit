//  Module: S_BOX
//
module S_BOX
    /*  package imports  */
    (
        input [31:0] word_in,  /*the row of matrix*/
        output [31:0] word_out
    );


    wire [7:0]S_MEM[0:255];


    assign word_out[31:24]=S_MEM[word_in[31:24]];
    assign word_out[23:16]=S_MEM[word_in[23:16]];
    assign word_out[15:8] =S_MEM[word_in[15:8]];
    assign word_out[7:0]  =S_MEM[word_in[7:0]];







    /*fill the memory table*/
  assign S_MEM[8'h00] = 8'h63;
  assign S_MEM[8'h01] = 8'h7c;
  assign S_MEM[8'h02] = 8'h77;
  assign S_MEM[8'h03] = 8'h7b;
  assign S_MEM[8'h04] = 8'hf2;
  assign S_MEM[8'h05] = 8'h6b;
  assign S_MEM[8'h06] = 8'h6f;
  assign S_MEM[8'h07] = 8'hc5;
  assign S_MEM[8'h08] = 8'h30;
  assign S_MEM[8'h09] = 8'h01;
  assign S_MEM[8'h0a] = 8'h67;
  assign S_MEM[8'h0b] = 8'h2b;
  assign S_MEM[8'h0c] = 8'hfe;
  assign S_MEM[8'h0d] = 8'hd7;
  assign S_MEM[8'h0e] = 8'hab;
  assign S_MEM[8'h0f] = 8'h76;
  assign S_MEM[8'h10] = 8'hca;
  assign S_MEM[8'h11] = 8'h82;
  assign S_MEM[8'h12] = 8'hc9;
  assign S_MEM[8'h13] = 8'h7d;
  assign S_MEM[8'h14] = 8'hfa;
  assign S_MEM[8'h15] = 8'h59;
  assign S_MEM[8'h16] = 8'h47;
  assign S_MEM[8'h17] = 8'hf0;
  assign S_MEM[8'h18] = 8'had;
  assign S_MEM[8'h19] = 8'hd4;
  assign S_MEM[8'h1a] = 8'ha2;
  assign S_MEM[8'h1b] = 8'haf;
  assign S_MEM[8'h1c] = 8'h9c;
  assign S_MEM[8'h1d] = 8'ha4;
  assign S_MEM[8'h1e] = 8'h72;
  assign S_MEM[8'h1f] = 8'hc0;
  assign S_MEM[8'h20] = 8'hb7;
  assign S_MEM[8'h21] = 8'hfd;
  assign S_MEM[8'h22] = 8'h93;
  assign S_MEM[8'h23] = 8'h26;
  assign S_MEM[8'h24] = 8'h36;
  assign S_MEM[8'h25] = 8'h3f;
  assign S_MEM[8'h26] = 8'hf7;
  assign S_MEM[8'h27] = 8'hcc;
  assign S_MEM[8'h28] = 8'h34;
  assign S_MEM[8'h29] = 8'ha5;
  assign S_MEM[8'h2a] = 8'he5;
  assign S_MEM[8'h2b] = 8'hf1;
  assign S_MEM[8'h2c] = 8'h71;
  assign S_MEM[8'h2d] = 8'hd8;
  assign S_MEM[8'h2e] = 8'h31;
  assign S_MEM[8'h2f] = 8'h15;
  assign S_MEM[8'h30] = 8'h04;
  assign S_MEM[8'h31] = 8'hc7;
  assign S_MEM[8'h32] = 8'h23;
  assign S_MEM[8'h33] = 8'hc3;
  assign S_MEM[8'h34] = 8'h18;
  assign S_MEM[8'h35] = 8'h96;
  assign S_MEM[8'h36] = 8'h05;
  assign S_MEM[8'h37] = 8'h9a;
  assign S_MEM[8'h38] = 8'h07;
  assign S_MEM[8'h39] = 8'h12;
  assign S_MEM[8'h3a] = 8'h80;
  assign S_MEM[8'h3b] = 8'he2;
  assign S_MEM[8'h3c] = 8'heb;
  assign S_MEM[8'h3d] = 8'h27;
  assign S_MEM[8'h3e] = 8'hb2;
  assign S_MEM[8'h3f] = 8'h75;
  assign S_MEM[8'h40] = 8'h09;
  assign S_MEM[8'h41] = 8'h83;
  assign S_MEM[8'h42] = 8'h2c;
  assign S_MEM[8'h43] = 8'h1a;
  assign S_MEM[8'h44] = 8'h1b;
  assign S_MEM[8'h45] = 8'h6e;
  assign S_MEM[8'h46] = 8'h5a;
  assign S_MEM[8'h47] = 8'ha0;
  assign S_MEM[8'h48] = 8'h52;
  assign S_MEM[8'h49] = 8'h3b;
  assign S_MEM[8'h4a] = 8'hd6;
  assign S_MEM[8'h4b] = 8'hb3;
  assign S_MEM[8'h4c] = 8'h29;
  assign S_MEM[8'h4d] = 8'he3;
  assign S_MEM[8'h4e] = 8'h2f;
  assign S_MEM[8'h4f] = 8'h84;
  assign S_MEM[8'h50] = 8'h53;
  assign S_MEM[8'h51] = 8'hd1;
  assign S_MEM[8'h52] = 8'h00;
  assign S_MEM[8'h53] = 8'hed;
  assign S_MEM[8'h54] = 8'h20;
  assign S_MEM[8'h55] = 8'hfc;
  assign S_MEM[8'h56] = 8'hb1;
  assign S_MEM[8'h57] = 8'h5b;
  assign S_MEM[8'h58] = 8'h6a;
  assign S_MEM[8'h59] = 8'hcb;
  assign S_MEM[8'h5a] = 8'hbe;
  assign S_MEM[8'h5b] = 8'h39;
  assign S_MEM[8'h5c] = 8'h4a;
  assign S_MEM[8'h5d] = 8'h4c;
  assign S_MEM[8'h5e] = 8'h58;
  assign S_MEM[8'h5f] = 8'hcf;
  assign S_MEM[8'h60] = 8'hd0;
  assign S_MEM[8'h61] = 8'hef;
  assign S_MEM[8'h62] = 8'haa;
  assign S_MEM[8'h63] = 8'hfb;
  assign S_MEM[8'h64] = 8'h43;
  assign S_MEM[8'h65] = 8'h4d;
  assign S_MEM[8'h66] = 8'h33;
  assign S_MEM[8'h67] = 8'h85;
  assign S_MEM[8'h68] = 8'h45;
  assign S_MEM[8'h69] = 8'hf9;
  assign S_MEM[8'h6a] = 8'h02;
  assign S_MEM[8'h6b] = 8'h7f;
  assign S_MEM[8'h6c] = 8'h50;
  assign S_MEM[8'h6d] = 8'h3c;
  assign S_MEM[8'h6e] = 8'h9f;
  assign S_MEM[8'h6f] = 8'ha8;
  assign S_MEM[8'h70] = 8'h51;
  assign S_MEM[8'h71] = 8'ha3;
  assign S_MEM[8'h72] = 8'h40;
  assign S_MEM[8'h73] = 8'h8f;
  assign S_MEM[8'h74] = 8'h92;
  assign S_MEM[8'h75] = 8'h9d;
  assign S_MEM[8'h76] = 8'h38;
  assign S_MEM[8'h77] = 8'hf5;
  assign S_MEM[8'h78] = 8'hbc;
  assign S_MEM[8'h79] = 8'hb6;
  assign S_MEM[8'h7a] = 8'hda;
  assign S_MEM[8'h7b] = 8'h21;
  assign S_MEM[8'h7c] = 8'h10;
  assign S_MEM[8'h7d] = 8'hff;
  assign S_MEM[8'h7e] = 8'hf3;
  assign S_MEM[8'h7f] = 8'hd2;
  assign S_MEM[8'h80] = 8'hcd;
  assign S_MEM[8'h81] = 8'h0c;
  assign S_MEM[8'h82] = 8'h13;
  assign S_MEM[8'h83] = 8'hec;
  assign S_MEM[8'h84] = 8'h5f;
  assign S_MEM[8'h85] = 8'h97;
  assign S_MEM[8'h86] = 8'h44;
  assign S_MEM[8'h87] = 8'h17;
  assign S_MEM[8'h88] = 8'hc4;
  assign S_MEM[8'h89] = 8'ha7;
  assign S_MEM[8'h8a] = 8'h7e;
  assign S_MEM[8'h8b] = 8'h3d;
  assign S_MEM[8'h8c] = 8'h64;
  assign S_MEM[8'h8d] = 8'h5d;
  assign S_MEM[8'h8e] = 8'h19;
  assign S_MEM[8'h8f] = 8'h73;
  assign S_MEM[8'h90] = 8'h60;
  assign S_MEM[8'h91] = 8'h81;
  assign S_MEM[8'h92] = 8'h4f;
  assign S_MEM[8'h93] = 8'hdc;
  assign S_MEM[8'h94] = 8'h22;
  assign S_MEM[8'h95] = 8'h2a;
  assign S_MEM[8'h96] = 8'h90;
  assign S_MEM[8'h97] = 8'h88;
  assign S_MEM[8'h98] = 8'h46;
  assign S_MEM[8'h99] = 8'hee;
  assign S_MEM[8'h9a] = 8'hb8;
  assign S_MEM[8'h9b] = 8'h14;
  assign S_MEM[8'h9c] = 8'hde;
  assign S_MEM[8'h9d] = 8'h5e;
  assign S_MEM[8'h9e] = 8'h0b;
  assign S_MEM[8'h9f] = 8'hdb;
  assign S_MEM[8'ha0] = 8'he0;
  assign S_MEM[8'ha1] = 8'h32;
  assign S_MEM[8'ha2] = 8'h3a;
  assign S_MEM[8'ha3] = 8'h0a;
  assign S_MEM[8'ha4] = 8'h49;
  assign S_MEM[8'ha5] = 8'h06;
  assign S_MEM[8'ha6] = 8'h24;
  assign S_MEM[8'ha7] = 8'h5c;
  assign S_MEM[8'ha8] = 8'hc2;
  assign S_MEM[8'ha9] = 8'hd3;
  assign S_MEM[8'haa] = 8'hac;
  assign S_MEM[8'hab] = 8'h62;
  assign S_MEM[8'hac] = 8'h91;
  assign S_MEM[8'had] = 8'h95;
  assign S_MEM[8'hae] = 8'he4;
  assign S_MEM[8'haf] = 8'h79;
  assign S_MEM[8'hb0] = 8'he7;
  assign S_MEM[8'hb1] = 8'hc8;
  assign S_MEM[8'hb2] = 8'h37;
  assign S_MEM[8'hb3] = 8'h6d;
  assign S_MEM[8'hb4] = 8'h8d;
  assign S_MEM[8'hb5] = 8'hd5;
  assign S_MEM[8'hb6] = 8'h4e;
  assign S_MEM[8'hb7] = 8'ha9;
  assign S_MEM[8'hb8] = 8'h6c;
  assign S_MEM[8'hb9] = 8'h56;
  assign S_MEM[8'hba] = 8'hf4;
  assign S_MEM[8'hbb] = 8'hea;
  assign S_MEM[8'hbc] = 8'h65;
  assign S_MEM[8'hbd] = 8'h7a;
  assign S_MEM[8'hbe] = 8'hae;
  assign S_MEM[8'hbf] = 8'h08;
  assign S_MEM[8'hc0] = 8'hba;
  assign S_MEM[8'hc1] = 8'h78;
  assign S_MEM[8'hc2] = 8'h25;
  assign S_MEM[8'hc3] = 8'h2e;
  assign S_MEM[8'hc4] = 8'h1c;
  assign S_MEM[8'hc5] = 8'ha6;
  assign S_MEM[8'hc6] = 8'hb4;
  assign S_MEM[8'hc7] = 8'hc6;
  assign S_MEM[8'hc8] = 8'he8;
  assign S_MEM[8'hc9] = 8'hdd;
  assign S_MEM[8'hca] = 8'h74;
  assign S_MEM[8'hcb] = 8'h1f;
  assign S_MEM[8'hcc] = 8'h4b;
  assign S_MEM[8'hcd] = 8'hbd;
  assign S_MEM[8'hce] = 8'h8b;
  assign S_MEM[8'hcf] = 8'h8a;
  assign S_MEM[8'hd0] = 8'h70;
  assign S_MEM[8'hd1] = 8'h3e;
  assign S_MEM[8'hd2] = 8'hb5;
  assign S_MEM[8'hd3] = 8'h66;
  assign S_MEM[8'hd4] = 8'h48;
  assign S_MEM[8'hd5] = 8'h03;
  assign S_MEM[8'hd6] = 8'hf6;
  assign S_MEM[8'hd7] = 8'h0e;
  assign S_MEM[8'hd8] = 8'h61;
  assign S_MEM[8'hd9] = 8'h35;
  assign S_MEM[8'hda] = 8'h57;
  assign S_MEM[8'hdb] = 8'hb9;
  assign S_MEM[8'hdc] = 8'h86;
  assign S_MEM[8'hdd] = 8'hc1;
  assign S_MEM[8'hde] = 8'h1d;
  assign S_MEM[8'hdf] = 8'h9e;
  assign S_MEM[8'he0] = 8'he1;
  assign S_MEM[8'he1] = 8'hf8;
  assign S_MEM[8'he2] = 8'h98;
  assign S_MEM[8'he3] = 8'h11;
  assign S_MEM[8'he4] = 8'h69;
  assign S_MEM[8'he5] = 8'hd9;
  assign S_MEM[8'he6] = 8'h8e;
  assign S_MEM[8'he7] = 8'h94;
  assign S_MEM[8'he8] = 8'h9b;
  assign S_MEM[8'he9] = 8'h1e;
  assign S_MEM[8'hea] = 8'h87;
  assign S_MEM[8'heb] = 8'he9;
  assign S_MEM[8'hec] = 8'hce;
  assign S_MEM[8'hed] = 8'h55;
  assign S_MEM[8'hee] = 8'h28;
  assign S_MEM[8'hef] = 8'hdf;
  assign S_MEM[8'hf0] = 8'h8c;
  assign S_MEM[8'hf1] = 8'ha1;
  assign S_MEM[8'hf2] = 8'h89;
  assign S_MEM[8'hf3] = 8'h0d;
  assign S_MEM[8'hf4] = 8'hbf;
  assign S_MEM[8'hf5] = 8'he6;
  assign S_MEM[8'hf6] = 8'h42;
  assign S_MEM[8'hf7] = 8'h68;
  assign S_MEM[8'hf8] = 8'h41;
  assign S_MEM[8'hf9] = 8'h99;
  assign S_MEM[8'hfa] = 8'h2d;
  assign S_MEM[8'hfb] = 8'h0f;
  assign S_MEM[8'hfc] = 8'hb0;
  assign S_MEM[8'hfd] = 8'h54;
  assign S_MEM[8'hfe] = 8'hbb;
  assign S_MEM[8'hff] = 8'h16;
    
endmodule: S_BOX
